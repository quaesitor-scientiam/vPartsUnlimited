module main

pub const module_name = 'main'
