module logging

pub const module_name = 'logging'
